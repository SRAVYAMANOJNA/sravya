    � B2SPICE zzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz    ��  CPart        S   �  ,      S   �  ,              Ammeter��  CIntPin    ��  CWire     �       �         �   @        �   @              BF469 �   �    	 �    
    �       �   �   �      �   �   �              resistor_generic �   �    �       4  �      �       S   �  ,      S   �  ,              Ammeter�    �     �       3  ��   CBehPin �  M+        R  M+����                        ��� �+  emitter      �	  emitter����                        �� 3    3  ��  CExtPin    ��  CVertex   @  �   ��  CSegment	   �   �  �   �   �   �  @                          �
    �   �  �   !                        �   M+x ��   �   �
  �   �   �   �
  `   �   & �   @  `   �   ( �   @   
   �   �   �   
   +        *     )         '         �   �   �
      -     &     %         $              �  �   M-��� @  �          VAm2    	 ��   CPin                   ��                                                           @   M+/�                   ��                                                      �   @   M-��  TLine �   @   �   @     ��                                                        2�     @       @     ��                                                        2� 4   X   `   X     ��                                                        �� 
 TRectangle        �   d                   ����                                                �   d   ��  TPolygon ����������������  ��          @ @                                           ��  TPointd   X        :�X   P    or  :�X   `        @ @ ��  
 TTextField $   $   �   L     ��                                                      $   $   �   L   $   $   �   L   [value]                       $   $   �   L   >�     �����        ��                                                           �����          �����      	[refname]       �  �  �	  <      �����       7   0 ? 1   5   @ 9 4   3 	     Ammeter     Miscellaneous      �?       ��   CAmmeterBehavior     ��  CValue ����    �i��       �������� M+M-  � �  M-      R  M-����                        ��AmmeterAmmeter   �             E Analog Meters   Generic   VAm2VAm2          ����  VAm ��   CPartPin    ����M+M+      PASAM+        F�   ����M-M-      PASAM-00E-   Analog MetersAmmeterGeneric              4  � �  M-      R  M-����                        ��E � �,  R-      
  R-����                        �� 4   4 �    �   �  �   �    �   �  �   M �   N �   �  �   O                 L                    �   R+    �   ,       @  R-    �  �         R1     /�                    ��                                                           @   R+/�                   ��                                                          �   R-2�     �   �����     ��    ��?                                                 2�    �   �����     ��    ��?                                                 2�    �   �����     ��    ��?                                                 2�    x   �����     ��                                                        2�    x   ����l     ��    `��                                                2�    `       X     ��    ��?                                                 2�     @       X     ��                                                        2�    `   ����l    	 ��        	                                                2�     �       �    
 ��        
                                                >�     t   �   �     ��                                                           t   �   �       t   �   �   [resistance]       @  <	  �  �	      `   �   �   >�     @   �   d     ��                                                           @   �   d       @   �   d   	[refname]       @  �  �  @	          t   $    R S T U V W X Y Z [ \ ] ^  �  resistor    resistor DINMiscellaneous      �?       ��  CResistorBehavior     C� ����     @�@1K      ��������C� ���� 27     ��������C� ����       ��������C� ����       �������� R+R- � �,  R+        
  R+����                        ��J resistorresistor                e J Passive   Generic   R1R1          ����    R F�    ����R+R+      PASAR+ 
G6    F�   ����R-R-      PASAR-(e�   Passive Generic              5  � �+  base      �	  base����                        ��e  5    5  �    P       �  Base    �   �   �  �   �   �
   �  `   l �   m �    @  `   n                  k               �   �  	Collector   �       �   @  Emitter    �             Q1     /�                   ��                                                           �   Base/�                   ��                                                      @   �   	Collector/�                    ��                                                      @   �   Emitter2�     �       �     ��                                                        2�     �       �     ��                                                        2�     �   0   �     ��    ��?                                                 2� @   �   0   �     ��                                                        2�     �   0   �     ��    ��?                                                 2� 0   �   @   �     ��                                                        2� 8   �   <   �    
 ��       	                                                2� 0   �   <   �     ��       
                                                >� .   H   �   h     ��                                                       .   H   �   h   .   H   �   h   
beta= [bf]       j  �  "  n      X   |   x   >� x      x       	 ��                                                      x      x      x      x              H    `  �  x      x      >�     4   x   X     ��                                                           4   x   X       4   x   X   	[refname]       �  �  h  <      4   x   X   >�        x   4     ��                                                              x   4          x   4   	[devname]        ����������������       x   4    s t u v w {   | x }   y   ~  z                 r   q      BJT npn     Miscellaneous      �?       ��  CBJTBehavior     C� ����        ��������C� ����       ��������C� ����       ��������C� ����       ��������C� ����       ��������C� ����  .     �������� 	collectorbaseemitter � �+  	collector        �	  	collector����                        ��h  �  �+  	substrate      �	  base����                        ��qbf469qbf469               � h  � 
Transistor1   Philips   Q1Q1                Q F�    ����	Collector	collector      PASAC( )    F�   ����Basebase      PASAB�e�   F�   ����Emitteremitter      PASAENDDA   F�   ����Base	substrate       PASABaseAM2.   
TransistorHigh Voltage NPN TransistorPhilipsTO-126             6  � �  M+        R  M+����                        ���  6    6  �    o        �   M+    �   &   �  �   M-    @  �          VAm1    	 /�                   ��                                                           @   M+/�                   ��                                                      �   @   M-2� �   @   �   @     ��    8��                                                2�     @       @     ��                                                        2� 4   X   `   X     ��    ��?                                                 6�        �   d                   ����                                                �   d   8� ����������������  ��          @ @                                           :�d   X        :�X   P    or  :�X   `        @ @ >� $   $   �   L     ��                                                      $   $   �   L   $   $   �   L   [value]                       $   $   �   L   >�     �����        ��                                                           �����          �����      	[refname]       �  |  �	        �����       �   � � �   �   � � �   � 	     Ammeter     Miscellaneous      �?       A�     C� ����    �i��       �������� M+M- � I AmmeterAmmeter   �            � I Analog Meters   Generic   VAm1VAm1          ����  VAm F�    ����M+M+      PASAM+@w�    F�   ����M-M-      PASAM-1.I    Analog MetersAmmeterGeneric                    �              
    M O l n       %   ! - ' ) +    o &  $ P k   , L   m N      " . ( *          ��  CLetter    6�  �  �  s      ����Arial����                       Arial     ��   4�  �	  �  3
      ����Arial����                       Arial     ��   3�    �  �      ����Arial����                       Arial     ��   50  0  �  �    �?����Arial����                       Arial            
 C�@ ����        ��������C�             0     ��������C� ����      @5     ��������C�  ʚ;�������?.1     ��������C�@ ����       ��������C� ����       ��������C� ����       ��������C� ����       ��������C� ���� true
     ��������C� ����  false     ��������               
                  C� ����        ��������C� ����       ��������C�  ����       ��������C�@ ����       ��������C�@ ����       ��������               
                  C� ����        ��������C� ����       ��������C�@ ����       ��������C�  ����       ��������C� ����       ��������C� ����       ��������C� ����       ��������C� ����       ��������C� ����       ��������C� ����       ��������C� ����       ��������               
                 C� ����dec     ��������C� ����     @�@1k     ��������C� ����    ��.A1meg     ��������C� ����       20     ��������C� ���� true     ��������C� ���� true     ��������C� ���� true	     ��������C� ����  false
     ��������               
                 C�  ����        ��������C�  ����       ��������C�  ����       ��������C� ����dec     ��������C� ����       ��������C� ����       ��������C� ����  	     ��������C� ����  
     ��������               
                  	 C� ����        ��������C� ����       ��������C� ����       ��������C� ����       ��������C� ����       ��������C� ����       ��������C� ����       ��������C� ����       ��������C� ����       ��������               
                 C� ����        ��������C� ����       ��������C� ����       ��������C� ����dec     ��������C� ����       ��������               
                    C�             0      ��������C� ��� ����MbP?1m     ��������C� �� �h㈵��>10u     ��������C� '  ���ư>1u     ��������C� ���� True     ��������C� ����  F     ��������C� ���� true     ��������C� ����  false     ��������               
                 C� ����     @�@1K      ��������C�  ����       ��������C�  ����       ��������C�  ����       ��������               
         ��              C�  ����        ��������              
                  C�  ����        ��������              
                                  
                 C�@ ����        ��������C�@ ����       ��������C� ����       ��������C� ����       ��������C� ����       ��������C� ����       ��������C� ����       ��������C� ����       ��������C� ����       ��������C� ���� true	     ��������C� ����  false
     ��������C� ���� true     ��������C� ����  false     ��������               
                 C� ����       5      ��������C� ����       5     ��������C� ����       5     ��������C� ����       5     ��������C� ����       ��������C� ����  	     ��������C� ����  
     ��������C� ����       ��������C� ����       ��������C� ����       ��������C� ���� true     ��������C�@ ����       ��������C�@ ����       ��������C� ����       ��������C� ����       ��������C� ����       ��������C� ����dec     ��������C� ����       ��������C� ����       ��������C� ����       ��������C� ���� true     ��������C� ���� true     ��������C� ���� true     ��������C� ����  false     ��������C� ���� true     ��������C� ����  false      ��������C� ���� true!     ��������C� ����  false"     ��������               
                        C� ����       5      ��������C� ����       5     ��������C� ����       5     ��������C� ����       5     ��������C� ����       ��������C� ����  	     ��������C� ����  
     ��������C� ����       ��������C� ����       ��������C� ����       ��������C� ���� true     ��������C�@ ����       ��������C�@ ����       ��������C� ����       ��������C� ����       ��������C� ����       ��������C� ����dec     ��������C� ����       ��������C� ����       ��������C� ����       ��������C� ���� true     ��������C� ���� true     ��������C� ���� true     ��������C� ����  false     ��������C� ���� true     ��������C� ����  false      ��������C� ���� true!     ��������C� ����  false"     ��������               
                 C� ����       5      ��������C� ����       5     ��������C� ����       5     ��������C� ����       5     ��������C� ����       ��������C� ����  	     ��������C� ����  
     ��������C� ����       ��������C� ����       ��������C� ����       ��������C� ���� true     ��������C�@ ����       ��������C�@ ����       ��������C� ����       ��������C� ����       ��������C� ����       ��������C� ����dec     ��������C� ����       ��������C� ����       ��������C� ����       ��������C� ���� true     ��������C� ���� true     ��������C� ���� true     ��������C� ����  false     ��������C� ���� true     ��������C� ����  false      ��������C� ���� true!     ��������C� ����  false"     ��������               
                 C� ����       5      ��������C� ����       5     ��������C� ����       5     ��������C� ����       5     ��������C� ����       ��������C� ����  	     ��������C� ����  
     ��������C� ����       ��������C� ����       ��������C� ����       ��������C� ���� true     ��������C�@ ����       ��������C�@ ����       ��������C� ����       ��������C� ����       ��������C� ����       ��������C� ����dec     ��������C� ����       ��������C� ����       ��������C� ����       ��������C� ���� true     ��������C� ���� true     ��������C� ���� true     ��������C� ����  false     ��������C� ���� true     ��������C� ����  false      ��������C� ���� true!     ��������C� ����  false"     ��������               
                 C�@ ����        ��������C�@ ����       ��������C� ����       ��������C� ����       ��������C� ����       ��������C� ����       ��������C� ����       ��������C� ����       ��������C� ����decade     ��������C� ���� true     ��������C� ���� true     ��������C� ���� true     ��������C� ����  false     ��������               
                 C� ����        ��������C� ����       ��������C�@ ����       ��������C�  ����       ��������C� ����       ��������C� ����       ��������C� ����       ��������C� ����       ��������C� ����       ��������C� ����       ��������C� ����       ��������               
                        C� ����dec     ��������C� ����     @�@1k     ��������C� ����    ��.A1meg     ��������C� ����       20     ��������C� ����        0     ��������C� ����        0     ��������C� ���� true	     ��������C� ���� true
     ��������C� ����      I@50     ��������C� ���� true     ��������C� ����  false     ��������               
                         / C� ���� x'     ��������C�     �-���q=1E-12     ��������C� @B -C��6?1E-4     ��������C� ���� x     ��������C� ���� x     ��������C� ���� x     ��������C� ���� x     ��������C� ���� x     ��������C� ���� x     ��������C� ���� x	     ��������C� ���� x!     ��������C� ����    �  500
     ��������C� ���� x     ��������C� ����    �  500     ��������C� ���� x$     ��������C� ���� x$     ��������C� ���� x%     ��������C� ���� x"     ��������C�  ���� x*     ��������C� ���� x     ��������C� ���� x     ��������C� ���� x     ��������C� ���� x&     ��������C� ���� x     ��������C� ���� x     ��������C� ���� x     ��������C� ���� x+     ��������C� ���� x,     ��������C� ���� x-     ��������C� ���� xg     ��������C� ���� xf     ��������C� ���� xd     ��������C� ���� xe     ��������C� ���� xh     ��������C� ���� xj     ��������C� ���� xi     ��������C� ���� xk     ��������C� ����    e��A1Gl     ��������C�             0�     ��������C� ����      @5�     ��������C� ����      @2.5�     ��������C� ����      �?.5�     ��������C� ����      @4.5�     ��������C� 
   ��&�.>1n�     ��������C� 
   ��&�.>1n�     ��������C� 
   ��&�.>1n�     ��������C� 
   ��&�.>1n�     ��������           ��  CPrimitiveModel    qbf469  , C� ���� t     ��������C� ����       ��������C�     ?۬���=	7.974e-15     ��������C� ����     �^@122     ��������C� ����-�����?0.993     ��������C� ������(\��9@25.51     ��������C�  !"4��k��?0.01029     ��������C�     L��>T�<	2.266e-16
     ��������C� �����z�G��?1.18     ��������C� ����q=
ף�@6.235     ��������C� ����+�����?0.999     ��������C� �����G�zn3@19.43     ��������C� @^u��gy�?0.02746     ��������C�     aM[�%�=4.33e-12     ��������C� ����'1�Z�?1.397     ��������C� ����      �?1     ��������C� '  ���ư>1e-06     ��������C� ����      �?0.5     ��������C� ����q���h�?0.3814     ��������C� ����j�t��?0.439     ��������C�     ז�IK'�=	1.742e-11     ��������C� ��������Q�?0.4581     ��������C� ����������?0.3092     ��������C�    ��zM>	7.073e-10     ��������C� ����     r@289.5     ��������C� �����~j�t�@6.144     ��������C� ��Y�A`��"�?0.1495      ��������C�             0!     ��������C�     8Oh?*0�=	5.045e-12"     ��������C� ��ku���K7�?0.197#     ��������C� ��t]�C����?0.1947%     ��������C� @f>J{�/L��?0.1041'     ��������C� d   :�0�yE>1e-08(     ��������C�             0)     ��������C�      0*     ��������C� ����      �?0.75+     ��������C� ����Zd;�O�?0.333-     ��������C�             0/     ��������C� ������(\���?1.110     ��������C� ����      @31     ��������C� �����K7�A`�?0.85552     ��������C� ���� 27;     ��������C�      0<     ��������C� ���� 1=     ��������    General Purpose NPN Transistor Philips��   CPrimitiveModelType &Junction Field effect transistor model����BJTQ>   ��  	 CParmDefn����  
NPN or PNP    Processtype         5    �����  NPN type device    Processnpn 0     e     �����  PNP type device    Processpnp 0     f     ����� 1.0e-16Saturation Current    ProcessisA0      g     ����� 100Ideal forward beta    Processbf 0      h     ����� 1.0Forward emission coefficient    Processnf 0      i     ����� infForward Early voltage    ProcessvafV0      j     ����� inf     ProcessvaV0     j     ����� inf$Forward beta roll-off corner current    ProcessikfA0      k     ����� inf     ProcessikA0    	 k     ����� 0B-E leakage saturation current    ProcessiseA0     
 l     ����� 1.5 B-E leakage emission coefficient    Processne 0      n     ����� 1Ideal reverse beta    Processbr 0      o     ����� 1Reverse emission coefficient    Processnr 0      p     ����� infReverse Early voltage    ProcessvarV0      q     ����� inf     ProcessvbV0     q     ����� inf$reverse beta roll-off corner current    ProcessikrA0      r     ����� 0B-C leakage saturation current    ProcessiscA0      s     ����� 2 B-C leakage emission coefficient    Processnc 0      u     ����� 0Zero bias base resistance    ProcessrbOhm0      v     ����� inf&Current for base resistance=(rb+rbm)/2    ProcessirbA0      w     ����� 0Minimum base resistance    ProcessrbmOhm0      x     ����� 0Emitter resistance    ProcessreOhm0      y     ����� 0Collector resistance    ProcessrcOhm0      z     ����� 0#Zero bias B-E depletion capacitance    ProcesscjeF0     {     ����� 0.75B-E built in potential    ProcessvjeV0     |     ����� 0.75     ProcesspeV0     |     ����� 0.33 B-E junction grading coefficient    Processmje 0     }     ����� 0.33     Processme 0     }     ����� 0Ideal forward transit time    Processtfsec0     ~     ����� 0%Coefficient for bias dependence of TF    Processxtf 0          ����� inf#Voltage giving VBC dependence of TF    ProcessvtfV0     �     ����� 0High current dependence of TF    ProcessitfA0      �     ����� 0Excess phase    Processptfdeg0    ! �     ����� 0#Zero bias B-C depletion capacitance    ProcesscjcF0    " �     ����� 0.75B-C built in potential    ProcessvjcV0    # �     �����       Processpc 0    $ �     ����� 0.33 B-C junction grading coefficient    Processmjc 0    % �     �����       Processmc 0    & �     ����� 1$Fraction of B-C cap to internal base    Processxcjc 0    ' �     ����� 0Ideal reverse transit time    Processtrsec0    ( �     ����� 0Zero bias C-S capacitance    ProcesscjsF0    ) �     ����� 0Zero bias C-S capacitance    ProcessccsF0    * �     ����� 0.75%Substrate junction built in potential    ProcessvjsV0    + �     ����� 0.75     ProcesspsV0    , �     ����� 0&Substrate junction grading coefficient    Processmjs 0    - �     ����� 0     Processms 0    . �     ����� 0#Forward and reverse beta temp. exp.    Processxtb 0     / �     ����� 1.11"Energy gap for IS temp. dependency    ProcessegeV0     0 �     ����� 3Temp. exponent for IS    Processxti 0     1 �     ����� 0.5#Forward bias junction fit parameter    Processfc 0     2 �     �����  Inverse early voltage:forward    Processinvearlyvoltf     3 -    �����  Inverse early voltage:reverse    Processinvearlyvoltr     4 .    �����  Inverse roll off - forward    Processinvrollofff     5 /    �����  Inverse roll off - reverse    Processinvrolloffr     6 0    �����  Collector conductance    Processcollectorconduct     7 1    �����  Emitter conductance    Processemitterconduct     8 2    �����  Transit time VBC factor    Processtranstimevbcfact     9 3    �����  Excess phase fact.    Processexcessphasefactor     : 4    ����� 27!Parameter measurement temperature    Processtnomdeg C0     ; �     ����� 0Flicker Noise Coefficient    Processkf 0     < �     ����� 1Flicker Noise Exponent    Processaf 0     = �        npnpnp��                      Ariald         �	     x� ��w           �	     x� ��w                        ����            ����                  ?             M�       ��  ?             M�       ��                ����                                  ?             M�        ��  ?             M�        ��                ����                                  ?             M�        ��  ?             M�        ��                ����                                  ?             M�        ��  ?             M�        ��                ����                                  ?             M�        ��  ?             M�        ��                ����                                  ?             M�        ��  ?             M�        ��                ����                                  ?             M�        ��  ?             M�        ��                ����                                  ?             M�        ��  ?             M�        ��                ����                                  ?             M�        ��  ?             M�        ��            	    ����                                  ?             M�        ��  ?             M�        ��            
    ����                                  ?             M�        ��  ?             M�        ��                ����                                  ?             M�        ��  ?             M�        ��                ����                                  ?             M�        ��  ?             M�        ��                ����                                  ?             M�        ��  ?             M�        ��                ����                                  ?             M�        ��  ?             M�        ��                ����                                  ?             M�        ��  ?             M�        ��                ����                                  ?             M�        ��  ?             M�        ��                ����                                  ?             M�        ��  ?             M�        ��                ����                                  ?             M�        ��  ?             M�        ��                ����                                  ?             M�        ��  ?             M�        ��                ����                                  ?             M�        ��  ?             M�        ��                ����                                  ?             M�        ��  ?             M�        ��                ����                                  ?             M�        ��  ?             M�        ��                ����                                  ?             M�        ��  ?             M�        ��                ����                                  ?             M�        ��  ?             M�        ��                ����                                  ?             M�        ��  ?             M�        ��                ����                                  ?             M�        ��  ?             M�        ��                ����                                  ?             M�        ��  ?             M�        ��                ����                                  ?             M�        ��  ?             M�        ��                ����                                 >          ��   CDigSimResTemplate                ���       ����  ����:�0�yU>20.00n���   ����                       Arial����                       Arial����                       Arial  �   �  �                                ����  ���� ������       ����  ���� ������                 �               ����  �����       200������         0.000000e+000��    ��������      0.000000e+000��    ��������      0.000000e+000��    ��������   ����                       Arial����                       Arial����                       Arial����                       Arial      �       �         �     �   �  �  Circuit1                  ����  ��    ��������                               3  TO-126�3 pin transistor package                                                                                                                                                                                                                                       ��   CPackageAliasSuperPCB TO-126    -�EagleNPN.LBRTO126    -�Orcad TO126    -�
UlitiboardUltilib.l55TO126    -�Eagletransistor-npnTO126    -�Eagletransistor-fetTO126    -�Eagletransistor-pnpTO126    -�Eagletransistor-powerTO126AV   ECB        A                      �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New� � �     �   �   �     �              H            �� H      $           H                           2         �  �                                      ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New� � �     �   �   �     �              H            �� H      $           H                           2         �  �                                      ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New� � �     �   �   �     �              H            �� H      $           H                           2         �  �                                      ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New� � �     �   �   �     �              H            �� H      $           H                           2         �  �                                      ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New� � �     �   �   �     �              H            �� H      $           H                           2         �  �                                      ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New� � �     �   �   �     �              H            �� H      $           H                           2         �  �                                      ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New� � �     �   �   �     �              H            �� H      $           H                           2         �  �                                      ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New� � �     �   �   �     �              H            �� H      $           H                           2         �  �                                      ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New� � �     �   �   �     �              H            �� H      $           H                           2         �  �                                      ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New� � �     �   �   �     �              H            �� H      $           H                           2         �  �                                      ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New� � �     �   �   �     �              H            �� H      $           H                           2         �  �                                      ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New� � �     �   �   �     �              H            �� H      $           H                           2         �  �                                      ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New� � �     �   �   �     �              H            �� H      $           H                           2         �  �                                      ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New� � �     �   �   �     �              H            �� H      $           H                           2         �  �                                      ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New� � �     �   �   �     �              H            �� H      $           H                           2         �  �                                      ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New� � �     �   �   �     �              H            �� H      $           H                           2         �  �                                      ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New� � �     �   �   �     �              H            �� H      $           H                           2         �  �                                      ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New� � �     �   �   �     �              H            �� H      $           H                           2         �  �                                      ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New� � �     �   �   �     �              H            �� H      $           H                           2         �  �                                      ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New� � �     �   �   �     �              H            �� H      $           H                           2         �  �                                      ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New� � �     �   �   �     �              H            �� H      $           H                           2         �  �                                      ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New� � �     �   �   �     �              H            �� H      $           H                           2         �  �                                      ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New� � �     �   �   �     �              H            �� H      $           H                           2         �  �                                      ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New� � �     �   �   �     �              H            �� H      $           H                           2         �  �                                      ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New� � �     �   �   �     �              H            �� H      $           H                           2         �  �                                      ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New� � �     �   �   �     �              H            �� H      $           H                           2         �  �                                      ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New� � �     �   �   �     �              H            �� H      $           H                           2         �  �                                      ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New� � �     �   �   �     �              H            �� H      $           H                           2         �  �                                      ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New� � �     �   �   �     �              H            �� H      $           H                           2         �  �                                      ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New� � �     �   �   �     �              H            �� H      $           H                           2         �  �                                      ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                               �� 	 CTitleBox                                                      �  �                6�         �  @                  ���                                                  �  @  2�     <   �  <     ��                                                        2�     |   �  |     ��                                                        2�     �   �  �     ��                                                        2�     �   �  �     ��                                                        >� �      �  4     ��                                                      �      �  4   �      �  4   [title]                                       >� �   D   �  t     ��                                                      �   D   �  t   �   D   �  t   [description]                                       >� `   �   h  �     ��                                                      `   �   h  �   `   �   h  �   [id]                                       >� �   �   �  �     ��                                                      �   �   �  �   �   �   �  �   
[designer]                                       >�      �   8    ��        	                                                   �   8       �   8  Date :       �    H
  �                  >� �     �  4   	 ��        
                                              �     �  4  �     �  4  [date]                                       >�       t   8    
 ��                                                            t   8         t   8   Title :       �    
  �                  >�    L   �   x     ��                                                         L   �   x      L   �   x   Description :       �  �  �  �                  >�    �   �   �     ��                                                         �   �   �      �   �   �   ID :       �  �  �	  P                  >�    �   �   �     ��                                                         �   �   �      �   �   �   
Designer :       �  \  8                     89:;<=>?@BCDEF          A     	title box    Analog Misc      �?    9 
 ��  CParamSubBehavior     C�  ����        ��������C�  ����       ��������C�  ����       ��������C�  ����       ��������C�  ����       ��������      
 9                                      ������   CParamSubModelType�� ����     �            title                �            description               �            id               �            designer               �            date                           ����            `         �?�� 	 CGraphDoc�  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New� � �     �   �   �     �                                                                                   2         �  �                                      ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                        �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New� � �     �   �   �     �                           D�vje     ATAB 1.0            03
LVAM1       ��  TSignal                      TIME� � � time                      W�                      i(vam1)� � � i(vam1)    TIME                 W�                      i(vam2)� �   i(vam2)    TIME                           2         �  �          Time                          ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                                                 